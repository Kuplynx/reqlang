module parser

import os
import net.http
/* Parses a req file into arguments for the client*/


pub fn parse_req(file_path string) ?http.FetchConfig {
	
}