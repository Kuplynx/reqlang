module parser

import regex
import http
import misc

/*
	The reqlang transpiler.
	Mostly using regular expressions, otto idc never said how I had to make it work, just be able to transpile the 
 */

fn create_var(line string) string {
	/*
		Creates a variable declaration from reqlang to V
		Regular variables are declared with 'mut', constants are not
		All types are inferred by the compiler, no need to specify
	 */
	if line.starts_with("const ") {
		return misc.convert_to_snake_case(line.replace("const ", "")).replace("=", ":=")
	} else {
		return "mut " + misc.convert_to_snake_case(line).replace("=", ":=")
	}
}

fn pass_one(code string) string {

	/*
		Pass one of the transpiler
		This section converts variables
	*/

	println("Pass 1, creating variables...")
	mut findvar_re, _, _ := regex.regex_base("([a-zA-Z0-9_]+) = \"([^\"]*)\";")
	mut transpiled := code.split("\n")
	for i, line in transpiled {
		if findvar_re.find_all_str(line) != [] {
			println("\u001b[32mFound variable assignment on line $i \u001b[0m")
			transpiled[i] = create_var(line)
		}
	}
	return transpiled.join("\n")

}

fn pass_two(code string) string {

	/*
		Pass two of the transpiler
		This section converts 'req' functions
	*/

	println("Pass 2, creating 'req' functions...")
	/* Some unnecessary steps have to be taken for it to work with V's regex engine, otherwise it will just segfault */
	mut findfunc_re, _, _ := regex.regex_base("req ([a-zA-Z0-9_]+)[\(]+([:= _a-zA-Z0-9]*)[\)]+ [\{]+([\n\t:=\"/._;a-zA-Z0-9 ]+)[\}]+")
	mut funcs := findfunc_re.find_all_str(code)
	for i in 0..funcs.len {
		println("\u001b[32mFound request function \u001b[0m")
		funcs[i] = http.translate(funcs[i].split("\n")).join("\n")

	}
	return funcs.join("\n")

}


pub fn transpile(code string) string{
	mut transpiled := pass_one(code)
	transpiled = pass_two(transpiled)
	return "/* Generated by reqlang */
module main

import net.http

$transpiled

	"
}